module JERICALLA (
	input [16:0] inst,
	output reg [31:0] out
);

endmodule